CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 230 30 200 9
-4 82 1288 688
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
-4 82 1288 688
211288082 384
0
6 Title:
5 Name:
0
0
0
10
9 Resistor~
219 297 324 0 1 5
0 0
0
0 0 864 0
2 1k
-7 -14 7 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8953 0 0
0
0
11 Signal Gen~
195 99 369 0 19 64
0 3 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1203982336 0 1065353216
20
1 100000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 832 0
5 -1/1V
-18 -30 17 -22
2 V1
-7 -40 7 -32
0
0
38 %D %1 %2 DC 0 SIN(0 1 100k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
4441 0 0
0
0
7 Ground~
168 135 423 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3618 0 0
0
0
10 Capacitor~
219 468 324 0 2 5
0 4 6
0
0 0 832 0
5 375nF
-17 -18 18 -10
2 C3
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6153 0 0
0
0
10 Capacitor~
219 360 324 0 2 5
0 5 4
0
0 0 832 0
6 3.33uF
-21 -18 21 -10
2 C2
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5394 0 0
0
0
10 Capacitor~
219 252 324 0 2 5
0 7 5
0
0 0 832 0
4 25uF
-14 -18 14 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7734 0 0
0
0
9 Resistor~
219 513 369 0 3 5
0 2 6 -1
0
0 0 864 90
2 1k
8 0 22 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9914 0 0
0
0
9 Resistor~
219 414 369 0 3 5
0 2 4 -1
0
0 0 864 90
2 1k
8 0 22 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3747 0 0
0
0
9 Resistor~
219 306 369 0 3 5
0 2 5 -1
0
0 0 864 90
2 1k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3549 0 0
0
0
9 Resistor~
219 180 324 0 2 5
0 3 7
0
0 0 864 0
2 1k
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7931 0 0
0
0
13
2 0 0 0 0 0 0 1 0 0 12 2
315 324
315 324
1 0 0 0 0 0 0 1 0 0 12 2
279 324
279 324
1 0 2 0 0 4096 0 3 0 0 6 3
135 417
135 416
134 416
1 0 2 0 0 12288 0 7 0 0 5 4
513 387
512 387
512 416
414 416
1 0 2 0 0 8192 0 8 0 0 6 3
414 387
414 416
305 416
2 1 2 0 0 12416 0 2 9 0 0 5
130 374
134 374
134 416
306 416
306 387
1 1 3 0 0 8320 0 10 2 0 0 4
162 324
134 324
134 364
130 364
2 0 4 0 0 4096 0 8 0 0 11 2
414 351
414 324
2 0 5 0 0 4096 0 9 0 0 12 2
306 351
306 324
2 2 6 0 0 8320 0 7 4 0 0 3
513 351
513 324
477 324
2 1 4 0 0 4224 0 5 4 0 0 2
369 324
459 324
1 2 5 0 0 4224 0 5 6 0 0 2
351 324
261 324
2 1 7 0 0 4224 0 10 6 0 0 2
198 324
243 324
0
0
8 0 0
0
0
0
0 0 0
0
0 0 0
100 1 1e-006 1e+009
0 5e-005 2e-007 2e-007
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
2228876 4290624 100 100 0 0
77 66 1457 786
0 71 1500 960
1454 66
77 66
1457 66
1457 786
0 0
6.49709e-315 4.43665e-315 0 1.62413e-314 6.50121e-315 6.50121e-315
12403 0
4 30 50
1
513 334
0 6 0 0 1	0 10 0 0
2360240 8419392 100 100 0 0
77 66 707 366
2 522 752 966
707 66
77 66
707 66
707 366
0 0
4.94359e-315 0 5.18397e-315 1.57939e-314 4.94359e-315 4.94359e-315
12409 0
4 0.001 0.5
1
513 329
0 6 0 0 1	0 10 0 0
919710 4290624 100 100 0 0
77 66 717 366
746 526 1496 970
707 66
77 66
707 66
707 366
0 0
5.53553e-315 4.85009e-315 0 1.62122e-314 5.53553e-315 5.53553e-315
12401 0
4 30 50
1
513 104
0 6 0 0 1	0 10 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
